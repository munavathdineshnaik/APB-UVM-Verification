baseseq
