apbenv
