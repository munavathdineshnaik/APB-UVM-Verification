basetest
