apbif
